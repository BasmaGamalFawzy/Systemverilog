// struct & union
