// blocking & non-blocking assignments


