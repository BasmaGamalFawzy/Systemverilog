// Create a 1D bit array of size 8.
// Initialize it with binary values. 
// Write a program that inverts each bit and displays both original and inverted values.
