//clocking block 